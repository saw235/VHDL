----------------------------------------------------------------------------------
-- Entity:        RAM
-- Written By:    Natalie Brock, Sarah Sternby, Saw Xue Zheng
-- Date Created:  2 Nov 2016
-- Description:   RAM with generic number of addresses with a generic bit width
--
-- Revision History (date, initials, description):
-- 	
--
-- Dependencies:
-------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity RAM is generic(n 			: integer := 8;
						    bit_width  : integer := 48;
							 bit_depth	: integer := 256);
    Port ( ADDRESS 	: in  STD_LOGIC_VECTOR(n-1 downto 0);
           DATA_in 	: in  STD_LOGIC_VECTOR(bit_width-1 downto 0);
           WE 		 	: in  STD_LOGIC;
			  RESET		: in  STD_LOGIC;
           CLK 		: in  STD_LOGIC;
           DATA_out  : out STD_LOGIC_VECTOR(bit_width-1 downto 0));
end RAM;

architecture Behavioral of RAM is
	type RAM_TYPE is ARRAY(0 to bit_depth-1) of STD_LOGIC_VECTOR(bit_width-1 downto 0);
	signal RAM : RAM_TYPE := ( x"000000000000",
										x"000000FFFFFF",
										x"000000FF0000",
										x"00000000FF00",
										x"0000000000FF",
										x"000000FFFF00",
										x"00000000FFFF",
										x"000000FF00FF",
										x"000000C0C0C0",
										x"000000808080",
										x"000000800000",
										x"000000808000",
										x"000000008000",
										x"000000800080",
										x"000000008080",
										x"000000000080",
										x"FFFFFF000000",
										x"FFFFFFFFFFFF",
										x"FFFFFFFF0000",
										x"FFFFFF00FF00",
										x"FFFFFF0000FF",
										x"FFFFFFFFFF00",
										x"FFFFFF00FFFF",
										x"FFFFFFFF00FF",
										x"FFFFFFC0C0C0",
										x"FFFFFF808080",
										x"FFFFFF800000",
										x"FFFFFF808000",
										x"FFFFFF008000",
										x"FFFFFF800080",
										x"FFFFFF008080",
										x"FFFFFF000080",
										x"FF0000000000",
										x"FF0000FFFFFF",
										x"FF0000FF0000",
										x"FF000000FF00",
										x"FF00000000FF",
										x"FF0000FFFF00",
										x"FF000000FFFF",
										x"FF0000FF00FF",
										x"FF0000C0C0C0",
										x"FF0000808080",
										x"FF0000800000",
										x"FF0000808000",
										x"FF0000008000",
										x"FF0000800080",
										x"FF0000008080",
										x"FF0000000080",
										x"00FF00000000",
										x"00FF00FFFFFF",
										x"00FF00FF0000",
										x"00FF0000FF00",
										x"00FF000000FF",
										x"00FF00FFFF00",
										x"00FF0000FFFF",
										x"00FF00FF00FF",
										x"00FF00C0C0C0",
										x"00FF00808080",
										x"00FF00800000",
										x"00FF00808000",
										x"00FF00008000",
										x"00FF00800080",
										x"00FF00008080",
										x"00FF00000080",
										x"0000FF000000",
										x"0000FFFFFFFF",
										x"0000FFFF0000",
										x"0000FF00FF00",
										x"0000FF0000FF",
										x"0000FFFFFF00",
										x"0000FF00FFFF",
										x"0000FFFF00FF",
										x"0000FFC0C0C0",
										x"0000FF808080",
										x"0000FF800000",
										x"0000FF808000",
										x"0000FF008000",
										x"0000FF800080",
										x"0000FF008080",
										x"0000FF000080",
										x"FFFF00000000",
										x"FFFF00FFFFFF",
										x"FFFF00FF0000",
										x"FFFF0000FF00",
										x"FFFF000000FF",
										x"FFFF00FFFF00",
										x"FFFF0000FFFF",
										x"FFFF00FF00FF",
										x"FFFF00C0C0C0",
										x"FFFF00808080",
										x"FFFF00800000",
										x"FFFF00808000",
										x"FFFF00008000",
										x"FFFF00800080",
										x"FFFF00008080",
										x"FFFF00000080",
										x"00FFFF000000",
										x"00FFFFFFFFFF",
										x"00FFFFFF0000",
										x"00FFFF00FF00",
										x"00FFFF0000FF",
										x"00FFFFFFFF00",
										x"00FFFF00FFFF",
										x"00FFFFFF00FF",
										x"00FFFFC0C0C0",
										x"00FFFF808080",
										x"00FFFF800000",
										x"00FFFF808000",
										x"00FFFF008000",
										x"00FFFF800080",
										x"00FFFF008080",
										x"00FFFF000080",
										x"FF00FF000000",
										x"FF00FFFFFFFF",
										x"FF00FFFF0000",
										x"FF00FF00FF00",
										x"FF00FF0000FF",
										x"FF00FFFFFF00",
										x"FF00FF00FFFF",
										x"FF00FFFF00FF",
										x"FF00FFC0C0C0",
										x"FF00FF808080",
										x"FF00FF800000",
										x"FF00FF808000",
										x"FF00FF008000",
										x"FF00FF800080",
										x"FF00FF008080",
										x"FF00FF000080",
										x"C0C0C0000000",
										x"C0C0C0FFFFFF",
										x"C0C0C0FF0000",
										x"C0C0C000FF00",
										x"C0C0C00000FF",
										x"C0C0C0FFFF00",
										x"C0C0C000FFFF",
										x"C0C0C0FF00FF",
										x"C0C0C0C0C0C0",
										x"C0C0C0808080",
										x"C0C0C0800000",
										x"C0C0C0808000",
										x"C0C0C0008000",
										x"C0C0C0800080",
										x"C0C0C0008080",
										x"C0C0C0000080",
										x"808080000000",
										x"808080FFFFFF",
										x"808080FF0000",
										x"80808000FF00",
										x"8080800000FF",
										x"808080FFFF00",
										x"80808000FFFF",
										x"808080FF00FF",
										x"808080C0C0C0",
										x"808080808080",
										x"808080800000",
										x"808080808000",
										x"808080008000",
										x"808080800080",
										x"808080008080",
										x"808080000080",
										x"800000000000",
										x"800000FFFFFF",
										x"800000FF0000",
										x"80000000FF00",
										x"8000000000FF",
										x"800000FFFF00",
										x"80000000FFFF",
										x"800000FF00FF",
										x"800000C0C0C0",
										x"800000808080",
										x"800000800000",
										x"800000808000",
										x"800000008000",
										x"800000800080",
										x"800000008080",
										x"800000000080",
										x"808000000000",
										x"808000FFFFFF",
										x"808000FF0000",
										x"80800000FF00",
										x"8080000000FF",
										x"808000FFFF00",
										x"80800000FFFF",
										x"808000FF00FF",
										x"808000C0C0C0",
										x"808000808080",
										x"808000800000",
										x"808000808000",
										x"808000008000",
										x"808000800080",
										x"808000008080",
										x"808000000080",
										x"008000000000",
										x"008000FFFFFF",
										x"008000FF0000",
										x"00800000FF00",
										x"0080000000FF",
										x"008000FFFF00",
										x"00800000FFFF",
										x"008000FF00FF",
										x"008000C0C0C0",
										x"008000808080",
										x"008000800000",
										x"008000808000",
										x"008000008000",
										x"008000800080",
										x"008000008080",
										x"008000000080",
										x"800080000000",
										x"800080FFFFFF",
										x"800080FF0000",
										x"80008000FF00",
										x"8000800000FF",
										x"800080FFFF00",
										x"80008000FFFF",
										x"800080FF00FF",
										x"800080C0C0C0",
										x"800080808080",
										x"800080800000",
										x"800080808000",
										x"800080008000",
										x"800080800080",
										x"800080008080",
										x"800080000080",
										x"008080000000",
										x"008080FFFFFF",
										x"008080FF0000",
										x"00808000FF00",
										x"0080800000FF",
										x"008080FFFF00",
										x"00808000FFFF",
										x"008080FF00FF",
										x"008080C0C0C0",
										x"008080808080",
										x"008080800000",
										x"008080808000",
										x"008080008000",
										x"008080800080",
										x"008080008080",
										x"008080000080",
										x"000080000000",
										x"000080FFFFFF",
										x"000080FF0000",
										x"00008000FF00",
										x"0000800000FF",
										x"000080FFFF00",
										x"00008000FFFF",
										x"000080FF00FF",
										x"000080C0C0C0",
										x"000080808080",
										x"000080800000",
										x"000080808000",
										x"000080008000",
										x"000080800080",
										x"000080008080",
										x"000080000080");
begin
	process (CLK) is
		begin
			if (CLK'event and (CLK = '1')) then
				if (WE='1') then
					RAM(to_integer(unsigned(ADDRESS))) <= DATA_in;
				end if;
				DATA_out <= RAM(to_integer(unsigned(ADDRESS)));
			end if;
	end process;


end Behavioral;

