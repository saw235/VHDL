----------------------------------------------------------------------------
-- Entity:        FindAverage_4bit_tb
-- Written By:    Saw Xue Zheng
-- Date Created:  9/10/2016
-- Description:   Testbench for FindAverage_4bit
--
-- Revision History (date, initials, description):
-- 	9 September 16, xps5001, file created.

-- Dependencies:
--		FindAverage_4bit
----------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY FindAverage_4bit_tb IS
END FindAverage_4bit_tb;
 
ARCHITECTURE behavior OF FindAverage_4bit_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT FindAverage_4bit
    PORT(
         A 			: IN  std_logic_vector(3 downto 0);
         B 			: IN  std_logic_vector(3 downto 0);
         C 			: IN  std_logic_vector(3 downto 0);
         D 			: IN  std_logic_vector(3 downto 0);
         AVERAGE 	: OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic_vector(3 downto 0) := (others => '0');
   signal B : std_logic_vector(3 downto 0) := (others => '0');
   signal C : std_logic_vector(3 downto 0) := (others => '0');
   signal D : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal AVERAGE : std_logic_vector(3 downto 0);



	type test_vector_type is array(0 to 624) of STD_LOGIC_VECTOR(19 downto 0);
	constant TEST_VECTOR : test_vector_type := (
   --A			B				C				D				AVERAGE
	"1000"	&	"1000"	&	"1000"	&	"1000"	&	"1000", -- Average = -8
	"1000"	&	"1000"	&	"1000"	&	"1001"	&	"1000", -- Average = -8
	"1000"	&	"1000"	&	"1000"	&	"0000"	&	"1010", -- Average = -6
	"1000"	&	"1000"	&	"1000"	&	"0001"	&	"1010", -- Average = -6
	"1000"	&	"1000"	&	"1000"	&	"0111"	&	"1100", -- Average = -4
	"1000"	&	"1000"	&	"1001"	&	"1000"	&	"1000", -- Average = -8
	"1000"	&	"1000"	&	"1001"	&	"1001"	&	"1000", -- Average = -8
	"1000"	&	"1000"	&	"1001"	&	"0000"	&	"1010", -- Average = -6
	"1000"	&	"1000"	&	"1001"	&	"0001"	&	"1010", -- Average = -6
	"1000"	&	"1000"	&	"1001"	&	"0111"	&	"1100", -- Average = -4
	"1000"	&	"1000"	&	"0000"	&	"1000"	&	"1010", -- Average = -6
	"1000"	&	"1000"	&	"0000"	&	"1001"	&	"1010", -- Average = -6
	"1000"	&	"1000"	&	"0000"	&	"0000"	&	"1100", -- Average = -4
	"1000"	&	"1000"	&	"0000"	&	"0001"	&	"1100", -- Average = -4
	"1000"	&	"1000"	&	"0000"	&	"0111"	&	"1110", -- Average = -2
	"1000"	&	"1000"	&	"0001"	&	"1000"	&	"1010", -- Average = -6
	"1000"	&	"1000"	&	"0001"	&	"1001"	&	"1010", -- Average = -6
	"1000"	&	"1000"	&	"0001"	&	"0000"	&	"1100", -- Average = -4
	"1000"	&	"1000"	&	"0001"	&	"0001"	&	"1100", -- Average = -4
	"1000"	&	"1000"	&	"0001"	&	"0111"	&	"1110", -- Average = -2
	"1000"	&	"1000"	&	"0111"	&	"1000"	&	"1100", -- Average = -4
	"1000"	&	"1000"	&	"0111"	&	"1001"	&	"1100", -- Average = -4
	"1000"	&	"1000"	&	"0111"	&	"0000"	&	"1110", -- Average = -2
	"1000"	&	"1000"	&	"0111"	&	"0001"	&	"1110", -- Average = -2
	"1000"	&	"1000"	&	"0111"	&	"0111"	&	"1111", -- Average = -1
	"1000"	&	"1001"	&	"1000"	&	"1000"	&	"1000", -- Average = -8
	"1000"	&	"1001"	&	"1000"	&	"1001"	&	"1000", -- Average = -8
	"1000"	&	"1001"	&	"1000"	&	"0000"	&	"1010", -- Average = -6
	"1000"	&	"1001"	&	"1000"	&	"0001"	&	"1010", -- Average = -6
	"1000"	&	"1001"	&	"1000"	&	"0111"	&	"1100", -- Average = -4
	"1000"	&	"1001"	&	"1001"	&	"1000"	&	"1000", -- Average = -8
	"1000"	&	"1001"	&	"1001"	&	"1001"	&	"1001", -- Average = -7
	"1000"	&	"1001"	&	"1001"	&	"0000"	&	"1010", -- Average = -6
	"1000"	&	"1001"	&	"1001"	&	"0001"	&	"1011", -- Average = -5
	"1000"	&	"1001"	&	"1001"	&	"0111"	&	"1100", -- Average = -4
	"1000"	&	"1001"	&	"0000"	&	"1000"	&	"1010", -- Average = -6
	"1000"	&	"1001"	&	"0000"	&	"1001"	&	"1010", -- Average = -6
	"1000"	&	"1001"	&	"0000"	&	"0000"	&	"1100", -- Average = -4
	"1000"	&	"1001"	&	"0000"	&	"0001"	&	"1100", -- Average = -4
	"1000"	&	"1001"	&	"0000"	&	"0111"	&	"1110", -- Average = -2
	"1000"	&	"1001"	&	"0001"	&	"1000"	&	"1010", -- Average = -6
	"1000"	&	"1001"	&	"0001"	&	"1001"	&	"1011", -- Average = -5
	"1000"	&	"1001"	&	"0001"	&	"0000"	&	"1100", -- Average = -4
	"1000"	&	"1001"	&	"0001"	&	"0001"	&	"1101", -- Average = -3
	"1000"	&	"1001"	&	"0001"	&	"0111"	&	"1110", -- Average = -2
	"1000"	&	"1001"	&	"0111"	&	"1000"	&	"1100", -- Average = -4
	"1000"	&	"1001"	&	"0111"	&	"1001"	&	"1100", -- Average = -4
	"1000"	&	"1001"	&	"0111"	&	"0000"	&	"1110", -- Average = -2
	"1000"	&	"1001"	&	"0111"	&	"0001"	&	"1110", -- Average = -2
	"1000"	&	"1001"	&	"0111"	&	"0111"	&	"0000", -- Average = 0
	"1000"	&	"0000"	&	"1000"	&	"1000"	&	"1010", -- Average = -6
	"1000"	&	"0000"	&	"1000"	&	"1001"	&	"1010", -- Average = -6
	"1000"	&	"0000"	&	"1000"	&	"0000"	&	"1100", -- Average = -4
	"1000"	&	"0000"	&	"1000"	&	"0001"	&	"1100", -- Average = -4
	"1000"	&	"0000"	&	"1000"	&	"0111"	&	"1110", -- Average = -2
	"1000"	&	"0000"	&	"1001"	&	"1000"	&	"1010", -- Average = -6
	"1000"	&	"0000"	&	"1001"	&	"1001"	&	"1010", -- Average = -6
	"1000"	&	"0000"	&	"1001"	&	"0000"	&	"1100", -- Average = -4
	"1000"	&	"0000"	&	"1001"	&	"0001"	&	"1100", -- Average = -4
	"1000"	&	"0000"	&	"1001"	&	"0111"	&	"1110", -- Average = -2
	"1000"	&	"0000"	&	"0000"	&	"1000"	&	"1100", -- Average = -4
	"1000"	&	"0000"	&	"0000"	&	"1001"	&	"1100", -- Average = -4
	"1000"	&	"0000"	&	"0000"	&	"0000"	&	"1110", -- Average = -2
	"1000"	&	"0000"	&	"0000"	&	"0001"	&	"1110", -- Average = -2
	"1000"	&	"0000"	&	"0000"	&	"0111"	&	"0000", -- Average = 0
	"1000"	&	"0000"	&	"0001"	&	"1000"	&	"1100", -- Average = -4
	"1000"	&	"0000"	&	"0001"	&	"1001"	&	"1100", -- Average = -4
	"1000"	&	"0000"	&	"0001"	&	"0000"	&	"1110", -- Average = -2
	"1000"	&	"0000"	&	"0001"	&	"0001"	&	"1110", -- Average = -2
	"1000"	&	"0000"	&	"0001"	&	"0111"	&	"0000", -- Average = 0
	"1000"	&	"0000"	&	"0111"	&	"1000"	&	"1110", -- Average = -2
	"1000"	&	"0000"	&	"0111"	&	"1001"	&	"1110", -- Average = -2
	"1000"	&	"0000"	&	"0111"	&	"0000"	&	"0000", -- Average = 0
	"1000"	&	"0000"	&	"0111"	&	"0001"	&	"0000", -- Average = 0
	"1000"	&	"0000"	&	"0111"	&	"0111"	&	"0010", -- Average = 2
	"1000"	&	"0001"	&	"1000"	&	"1000"	&	"1010", -- Average = -6
	"1000"	&	"0001"	&	"1000"	&	"1001"	&	"1010", -- Average = -6
	"1000"	&	"0001"	&	"1000"	&	"0000"	&	"1100", -- Average = -4
	"1000"	&	"0001"	&	"1000"	&	"0001"	&	"1100", -- Average = -4
	"1000"	&	"0001"	&	"1000"	&	"0111"	&	"1110", -- Average = -2
	"1000"	&	"0001"	&	"1001"	&	"1000"	&	"1010", -- Average = -6
	"1000"	&	"0001"	&	"1001"	&	"1001"	&	"1011", -- Average = -5
	"1000"	&	"0001"	&	"1001"	&	"0000"	&	"1100", -- Average = -4
	"1000"	&	"0001"	&	"1001"	&	"0001"	&	"1101", -- Average = -3
	"1000"	&	"0001"	&	"1001"	&	"0111"	&	"1110", -- Average = -2
	"1000"	&	"0001"	&	"0000"	&	"1000"	&	"1100", -- Average = -4
	"1000"	&	"0001"	&	"0000"	&	"1001"	&	"1100", -- Average = -4
	"1000"	&	"0001"	&	"0000"	&	"0000"	&	"1110", -- Average = -2
	"1000"	&	"0001"	&	"0000"	&	"0001"	&	"1110", -- Average = -2
	"1000"	&	"0001"	&	"0000"	&	"0111"	&	"0000", -- Average = 0
	"1000"	&	"0001"	&	"0001"	&	"1000"	&	"1100", -- Average = -4
	"1000"	&	"0001"	&	"0001"	&	"1001"	&	"1101", -- Average = -3
	"1000"	&	"0001"	&	"0001"	&	"0000"	&	"1110", -- Average = -2
	"1000"	&	"0001"	&	"0001"	&	"0001"	&	"1111", -- Average = -1
	"1000"	&	"0001"	&	"0001"	&	"0111"	&	"0000", -- Average = 0
	"1000"	&	"0001"	&	"0111"	&	"1000"	&	"1110", -- Average = -2
	"1000"	&	"0001"	&	"0111"	&	"1001"	&	"1110", -- Average = -2
	"1000"	&	"0001"	&	"0111"	&	"0000"	&	"0000", -- Average = 0
	"1000"	&	"0001"	&	"0111"	&	"0001"	&	"0000", -- Average = 0
	"1000"	&	"0001"	&	"0111"	&	"0111"	&	"0010", -- Average = 2
	"1000"	&	"0111"	&	"1000"	&	"1000"	&	"1100", -- Average = -4
	"1000"	&	"0111"	&	"1000"	&	"1001"	&	"1100", -- Average = -4
	"1000"	&	"0111"	&	"1000"	&	"0000"	&	"1110", -- Average = -2
	"1000"	&	"0111"	&	"1000"	&	"0001"	&	"1110", -- Average = -2
	"1000"	&	"0111"	&	"1000"	&	"0111"	&	"1111", -- Average = -1
	"1000"	&	"0111"	&	"1001"	&	"1000"	&	"1100", -- Average = -4
	"1000"	&	"0111"	&	"1001"	&	"1001"	&	"1100", -- Average = -4
	"1000"	&	"0111"	&	"1001"	&	"0000"	&	"1110", -- Average = -2
	"1000"	&	"0111"	&	"1001"	&	"0001"	&	"1110", -- Average = -2
	"1000"	&	"0111"	&	"1001"	&	"0111"	&	"0000", -- Average = 0
	"1000"	&	"0111"	&	"0000"	&	"1000"	&	"1110", -- Average = -2
	"1000"	&	"0111"	&	"0000"	&	"1001"	&	"1110", -- Average = -2
	"1000"	&	"0111"	&	"0000"	&	"0000"	&	"0000", -- Average = 0
	"1000"	&	"0111"	&	"0000"	&	"0001"	&	"0000", -- Average = 0
	"1000"	&	"0111"	&	"0000"	&	"0111"	&	"0010", -- Average = 2
	"1000"	&	"0111"	&	"0001"	&	"1000"	&	"1110", -- Average = -2
	"1000"	&	"0111"	&	"0001"	&	"1001"	&	"1110", -- Average = -2
	"1000"	&	"0111"	&	"0001"	&	"0000"	&	"0000", -- Average = 0
	"1000"	&	"0111"	&	"0001"	&	"0001"	&	"0000", -- Average = 0
	"1000"	&	"0111"	&	"0001"	&	"0111"	&	"0010", -- Average = 2
	"1000"	&	"0111"	&	"0111"	&	"1000"	&	"1111", -- Average = -1
	"1000"	&	"0111"	&	"0111"	&	"1001"	&	"0000", -- Average = 0
	"1000"	&	"0111"	&	"0111"	&	"0000"	&	"0010", -- Average = 2
	"1000"	&	"0111"	&	"0111"	&	"0001"	&	"0010", -- Average = 2
	"1000"	&	"0111"	&	"0111"	&	"0111"	&	"0011", -- Average = 3
	"1001"	&	"1000"	&	"1000"	&	"1000"	&	"1000", -- Average = -8
	"1001"	&	"1000"	&	"1000"	&	"1001"	&	"1000", -- Average = -8
	"1001"	&	"1000"	&	"1000"	&	"0000"	&	"1010", -- Average = -6
	"1001"	&	"1000"	&	"1000"	&	"0001"	&	"1010", -- Average = -6
	"1001"	&	"1000"	&	"1000"	&	"0111"	&	"1100", -- Average = -4
	"1001"	&	"1000"	&	"1001"	&	"1000"	&	"1000", -- Average = -8
	"1001"	&	"1000"	&	"1001"	&	"1001"	&	"1001", -- Average = -7
	"1001"	&	"1000"	&	"1001"	&	"0000"	&	"1010", -- Average = -6
	"1001"	&	"1000"	&	"1001"	&	"0001"	&	"1011", -- Average = -5
	"1001"	&	"1000"	&	"1001"	&	"0111"	&	"1100", -- Average = -4
	"1001"	&	"1000"	&	"0000"	&	"1000"	&	"1010", -- Average = -6
	"1001"	&	"1000"	&	"0000"	&	"1001"	&	"1010", -- Average = -6
	"1001"	&	"1000"	&	"0000"	&	"0000"	&	"1100", -- Average = -4
	"1001"	&	"1000"	&	"0000"	&	"0001"	&	"1100", -- Average = -4
	"1001"	&	"1000"	&	"0000"	&	"0111"	&	"1110", -- Average = -2
	"1001"	&	"1000"	&	"0001"	&	"1000"	&	"1010", -- Average = -6
	"1001"	&	"1000"	&	"0001"	&	"1001"	&	"1011", -- Average = -5
	"1001"	&	"1000"	&	"0001"	&	"0000"	&	"1100", -- Average = -4
	"1001"	&	"1000"	&	"0001"	&	"0001"	&	"1101", -- Average = -3
	"1001"	&	"1000"	&	"0001"	&	"0111"	&	"1110", -- Average = -2
	"1001"	&	"1000"	&	"0111"	&	"1000"	&	"1100", -- Average = -4
	"1001"	&	"1000"	&	"0111"	&	"1001"	&	"1100", -- Average = -4
	"1001"	&	"1000"	&	"0111"	&	"0000"	&	"1110", -- Average = -2
	"1001"	&	"1000"	&	"0111"	&	"0001"	&	"1110", -- Average = -2
	"1001"	&	"1000"	&	"0111"	&	"0111"	&	"0000", -- Average = 0
	"1001"	&	"1001"	&	"1000"	&	"1000"	&	"1000", -- Average = -8
	"1001"	&	"1001"	&	"1000"	&	"1001"	&	"1001", -- Average = -7
	"1001"	&	"1001"	&	"1000"	&	"0000"	&	"1010", -- Average = -6
	"1001"	&	"1001"	&	"1000"	&	"0001"	&	"1011", -- Average = -5
	"1001"	&	"1001"	&	"1000"	&	"0111"	&	"1100", -- Average = -4
	"1001"	&	"1001"	&	"1001"	&	"1000"	&	"1001", -- Average = -7
	"1001"	&	"1001"	&	"1001"	&	"1001"	&	"1001", -- Average = -7
	"1001"	&	"1001"	&	"1001"	&	"0000"	&	"1011", -- Average = -5
	"1001"	&	"1001"	&	"1001"	&	"0001"	&	"1011", -- Average = -5
	"1001"	&	"1001"	&	"1001"	&	"0111"	&	"1100", -- Average = -4
	"1001"	&	"1001"	&	"0000"	&	"1000"	&	"1010", -- Average = -6
	"1001"	&	"1001"	&	"0000"	&	"1001"	&	"1011", -- Average = -5
	"1001"	&	"1001"	&	"0000"	&	"0000"	&	"1100", -- Average = -4
	"1001"	&	"1001"	&	"0000"	&	"0001"	&	"1101", -- Average = -3
	"1001"	&	"1001"	&	"0000"	&	"0111"	&	"1110", -- Average = -2
	"1001"	&	"1001"	&	"0001"	&	"1000"	&	"1011", -- Average = -5
	"1001"	&	"1001"	&	"0001"	&	"1001"	&	"1011", -- Average = -5
	"1001"	&	"1001"	&	"0001"	&	"0000"	&	"1101", -- Average = -3
	"1001"	&	"1001"	&	"0001"	&	"0001"	&	"1101", -- Average = -3
	"1001"	&	"1001"	&	"0001"	&	"0111"	&	"1110", -- Average = -2
	"1001"	&	"1001"	&	"0111"	&	"1000"	&	"1100", -- Average = -4
	"1001"	&	"1001"	&	"0111"	&	"1001"	&	"1100", -- Average = -4
	"1001"	&	"1001"	&	"0111"	&	"0000"	&	"1110", -- Average = -2
	"1001"	&	"1001"	&	"0111"	&	"0001"	&	"1110", -- Average = -2
	"1001"	&	"1001"	&	"0111"	&	"0111"	&	"0000", -- Average = 0
	"1001"	&	"0000"	&	"1000"	&	"1000"	&	"1010", -- Average = -6
	"1001"	&	"0000"	&	"1000"	&	"1001"	&	"1010", -- Average = -6
	"1001"	&	"0000"	&	"1000"	&	"0000"	&	"1100", -- Average = -4
	"1001"	&	"0000"	&	"1000"	&	"0001"	&	"1100", -- Average = -4
	"1001"	&	"0000"	&	"1000"	&	"0111"	&	"1110", -- Average = -2
	"1001"	&	"0000"	&	"1001"	&	"1000"	&	"1010", -- Average = -6
	"1001"	&	"0000"	&	"1001"	&	"1001"	&	"1011", -- Average = -5
	"1001"	&	"0000"	&	"1001"	&	"0000"	&	"1100", -- Average = -4
	"1001"	&	"0000"	&	"1001"	&	"0001"	&	"1101", -- Average = -3
	"1001"	&	"0000"	&	"1001"	&	"0111"	&	"1110", -- Average = -2
	"1001"	&	"0000"	&	"0000"	&	"1000"	&	"1100", -- Average = -4
	"1001"	&	"0000"	&	"0000"	&	"1001"	&	"1100", -- Average = -4
	"1001"	&	"0000"	&	"0000"	&	"0000"	&	"1110", -- Average = -2
	"1001"	&	"0000"	&	"0000"	&	"0001"	&	"1110", -- Average = -2
	"1001"	&	"0000"	&	"0000"	&	"0111"	&	"0000", -- Average = 0
	"1001"	&	"0000"	&	"0001"	&	"1000"	&	"1100", -- Average = -4
	"1001"	&	"0000"	&	"0001"	&	"1001"	&	"1101", -- Average = -3
	"1001"	&	"0000"	&	"0001"	&	"0000"	&	"1110", -- Average = -2
	"1001"	&	"0000"	&	"0001"	&	"0001"	&	"1111", -- Average = -1
	"1001"	&	"0000"	&	"0001"	&	"0111"	&	"0000", -- Average = 0
	"1001"	&	"0000"	&	"0111"	&	"1000"	&	"1110", -- Average = -2
	"1001"	&	"0000"	&	"0111"	&	"1001"	&	"1110", -- Average = -2
	"1001"	&	"0000"	&	"0111"	&	"0000"	&	"0000", -- Average = 0
	"1001"	&	"0000"	&	"0111"	&	"0001"	&	"0000", -- Average = 0
	"1001"	&	"0000"	&	"0111"	&	"0111"	&	"0010", -- Average = 2
	"1001"	&	"0001"	&	"1000"	&	"1000"	&	"1010", -- Average = -6
	"1001"	&	"0001"	&	"1000"	&	"1001"	&	"1011", -- Average = -5
	"1001"	&	"0001"	&	"1000"	&	"0000"	&	"1100", -- Average = -4
	"1001"	&	"0001"	&	"1000"	&	"0001"	&	"1101", -- Average = -3
	"1001"	&	"0001"	&	"1000"	&	"0111"	&	"1110", -- Average = -2
	"1001"	&	"0001"	&	"1001"	&	"1000"	&	"1011", -- Average = -5
	"1001"	&	"0001"	&	"1001"	&	"1001"	&	"1011", -- Average = -5
	"1001"	&	"0001"	&	"1001"	&	"0000"	&	"1101", -- Average = -3
	"1001"	&	"0001"	&	"1001"	&	"0001"	&	"1101", -- Average = -3
	"1001"	&	"0001"	&	"1001"	&	"0111"	&	"1110", -- Average = -2
	"1001"	&	"0001"	&	"0000"	&	"1000"	&	"1100", -- Average = -4
	"1001"	&	"0001"	&	"0000"	&	"1001"	&	"1101", -- Average = -3
	"1001"	&	"0001"	&	"0000"	&	"0000"	&	"1110", -- Average = -2
	"1001"	&	"0001"	&	"0000"	&	"0001"	&	"1111", -- Average = -1
	"1001"	&	"0001"	&	"0000"	&	"0111"	&	"0000", -- Average = 0
	"1001"	&	"0001"	&	"0001"	&	"1000"	&	"1101", -- Average = -3
	"1001"	&	"0001"	&	"0001"	&	"1001"	&	"1101", -- Average = -3
	"1001"	&	"0001"	&	"0001"	&	"0000"	&	"1111", -- Average = -1
	"1001"	&	"0001"	&	"0001"	&	"0001"	&	"1111", -- Average = -1
	"1001"	&	"0001"	&	"0001"	&	"0111"	&	"0001", -- Average = 1
	"1001"	&	"0001"	&	"0111"	&	"1000"	&	"1110", -- Average = -2
	"1001"	&	"0001"	&	"0111"	&	"1001"	&	"1110", -- Average = -2
	"1001"	&	"0001"	&	"0111"	&	"0000"	&	"0000", -- Average = 0
	"1001"	&	"0001"	&	"0111"	&	"0001"	&	"0001", -- Average = 1
	"1001"	&	"0001"	&	"0111"	&	"0111"	&	"0010", -- Average = 2
	"1001"	&	"0111"	&	"1000"	&	"1000"	&	"1100", -- Average = -4
	"1001"	&	"0111"	&	"1000"	&	"1001"	&	"1100", -- Average = -4
	"1001"	&	"0111"	&	"1000"	&	"0000"	&	"1110", -- Average = -2
	"1001"	&	"0111"	&	"1000"	&	"0001"	&	"1110", -- Average = -2
	"1001"	&	"0111"	&	"1000"	&	"0111"	&	"0000", -- Average = 0
	"1001"	&	"0111"	&	"1001"	&	"1000"	&	"1100", -- Average = -4
	"1001"	&	"0111"	&	"1001"	&	"1001"	&	"1100", -- Average = -4
	"1001"	&	"0111"	&	"1001"	&	"0000"	&	"1110", -- Average = -2
	"1001"	&	"0111"	&	"1001"	&	"0001"	&	"1110", -- Average = -2
	"1001"	&	"0111"	&	"1001"	&	"0111"	&	"0000", -- Average = 0
	"1001"	&	"0111"	&	"0000"	&	"1000"	&	"1110", -- Average = -2
	"1001"	&	"0111"	&	"0000"	&	"1001"	&	"1110", -- Average = -2
	"1001"	&	"0111"	&	"0000"	&	"0000"	&	"0000", -- Average = 0
	"1001"	&	"0111"	&	"0000"	&	"0001"	&	"0000", -- Average = 0
	"1001"	&	"0111"	&	"0000"	&	"0111"	&	"0010", -- Average = 2
	"1001"	&	"0111"	&	"0001"	&	"1000"	&	"1110", -- Average = -2
	"1001"	&	"0111"	&	"0001"	&	"1001"	&	"1110", -- Average = -2
	"1001"	&	"0111"	&	"0001"	&	"0000"	&	"0000", -- Average = 0
	"1001"	&	"0111"	&	"0001"	&	"0001"	&	"0001", -- Average = 1
	"1001"	&	"0111"	&	"0001"	&	"0111"	&	"0010", -- Average = 2
	"1001"	&	"0111"	&	"0111"	&	"1000"	&	"0000", -- Average = 0
	"1001"	&	"0111"	&	"0111"	&	"1001"	&	"0000", -- Average = 0
	"1001"	&	"0111"	&	"0111"	&	"0000"	&	"0010", -- Average = 2
	"1001"	&	"0111"	&	"0111"	&	"0001"	&	"0010", -- Average = 2
	"1001"	&	"0111"	&	"0111"	&	"0111"	&	"0100", -- Average = 4
	"0000"	&	"1000"	&	"1000"	&	"1000"	&	"1010", -- Average = -6
	"0000"	&	"1000"	&	"1000"	&	"1001"	&	"1010", -- Average = -6
	"0000"	&	"1000"	&	"1000"	&	"0000"	&	"1100", -- Average = -4
	"0000"	&	"1000"	&	"1000"	&	"0001"	&	"1100", -- Average = -4
	"0000"	&	"1000"	&	"1000"	&	"0111"	&	"1110", -- Average = -2
	"0000"	&	"1000"	&	"1001"	&	"1000"	&	"1010", -- Average = -6
	"0000"	&	"1000"	&	"1001"	&	"1001"	&	"1010", -- Average = -6
	"0000"	&	"1000"	&	"1001"	&	"0000"	&	"1100", -- Average = -4
	"0000"	&	"1000"	&	"1001"	&	"0001"	&	"1100", -- Average = -4
	"0000"	&	"1000"	&	"1001"	&	"0111"	&	"1110", -- Average = -2
	"0000"	&	"1000"	&	"0000"	&	"1000"	&	"1100", -- Average = -4
	"0000"	&	"1000"	&	"0000"	&	"1001"	&	"1100", -- Average = -4
	"0000"	&	"1000"	&	"0000"	&	"0000"	&	"1110", -- Average = -2
	"0000"	&	"1000"	&	"0000"	&	"0001"	&	"1110", -- Average = -2
	"0000"	&	"1000"	&	"0000"	&	"0111"	&	"0000", -- Average = 0
	"0000"	&	"1000"	&	"0001"	&	"1000"	&	"1100", -- Average = -4
	"0000"	&	"1000"	&	"0001"	&	"1001"	&	"1100", -- Average = -4
	"0000"	&	"1000"	&	"0001"	&	"0000"	&	"1110", -- Average = -2
	"0000"	&	"1000"	&	"0001"	&	"0001"	&	"1110", -- Average = -2
	"0000"	&	"1000"	&	"0001"	&	"0111"	&	"0000", -- Average = 0
	"0000"	&	"1000"	&	"0111"	&	"1000"	&	"1110", -- Average = -2
	"0000"	&	"1000"	&	"0111"	&	"1001"	&	"1110", -- Average = -2
	"0000"	&	"1000"	&	"0111"	&	"0000"	&	"0000", -- Average = 0
	"0000"	&	"1000"	&	"0111"	&	"0001"	&	"0000", -- Average = 0
	"0000"	&	"1000"	&	"0111"	&	"0111"	&	"0010", -- Average = 2
	"0000"	&	"1001"	&	"1000"	&	"1000"	&	"1010", -- Average = -6
	"0000"	&	"1001"	&	"1000"	&	"1001"	&	"1010", -- Average = -6
	"0000"	&	"1001"	&	"1000"	&	"0000"	&	"1100", -- Average = -4
	"0000"	&	"1001"	&	"1000"	&	"0001"	&	"1100", -- Average = -4
	"0000"	&	"1001"	&	"1000"	&	"0111"	&	"1110", -- Average = -2
	"0000"	&	"1001"	&	"1001"	&	"1000"	&	"1010", -- Average = -6
	"0000"	&	"1001"	&	"1001"	&	"1001"	&	"1011", -- Average = -5
	"0000"	&	"1001"	&	"1001"	&	"0000"	&	"1100", -- Average = -4
	"0000"	&	"1001"	&	"1001"	&	"0001"	&	"1101", -- Average = -3
	"0000"	&	"1001"	&	"1001"	&	"0111"	&	"1110", -- Average = -2
	"0000"	&	"1001"	&	"0000"	&	"1000"	&	"1100", -- Average = -4
	"0000"	&	"1001"	&	"0000"	&	"1001"	&	"1100", -- Average = -4
	"0000"	&	"1001"	&	"0000"	&	"0000"	&	"1110", -- Average = -2
	"0000"	&	"1001"	&	"0000"	&	"0001"	&	"1110", -- Average = -2
	"0000"	&	"1001"	&	"0000"	&	"0111"	&	"0000", -- Average = 0
	"0000"	&	"1001"	&	"0001"	&	"1000"	&	"1100", -- Average = -4
	"0000"	&	"1001"	&	"0001"	&	"1001"	&	"1101", -- Average = -3
	"0000"	&	"1001"	&	"0001"	&	"0000"	&	"1110", -- Average = -2
	"0000"	&	"1001"	&	"0001"	&	"0001"	&	"1111", -- Average = -1
	"0000"	&	"1001"	&	"0001"	&	"0111"	&	"0000", -- Average = 0
	"0000"	&	"1001"	&	"0111"	&	"1000"	&	"1110", -- Average = -2
	"0000"	&	"1001"	&	"0111"	&	"1001"	&	"1110", -- Average = -2
	"0000"	&	"1001"	&	"0111"	&	"0000"	&	"0000", -- Average = 0
	"0000"	&	"1001"	&	"0111"	&	"0001"	&	"0000", -- Average = 0
	"0000"	&	"1001"	&	"0111"	&	"0111"	&	"0010", -- Average = 2
	"0000"	&	"0000"	&	"1000"	&	"1000"	&	"1100", -- Average = -4
	"0000"	&	"0000"	&	"1000"	&	"1001"	&	"1100", -- Average = -4
	"0000"	&	"0000"	&	"1000"	&	"0000"	&	"1110", -- Average = -2
	"0000"	&	"0000"	&	"1000"	&	"0001"	&	"1110", -- Average = -2
	"0000"	&	"0000"	&	"1000"	&	"0111"	&	"0000", -- Average = 0
	"0000"	&	"0000"	&	"1001"	&	"1000"	&	"1100", -- Average = -4
	"0000"	&	"0000"	&	"1001"	&	"1001"	&	"1100", -- Average = -4
	"0000"	&	"0000"	&	"1001"	&	"0000"	&	"1110", -- Average = -2
	"0000"	&	"0000"	&	"1001"	&	"0001"	&	"1110", -- Average = -2
	"0000"	&	"0000"	&	"1001"	&	"0111"	&	"0000", -- Average = 0
	"0000"	&	"0000"	&	"0000"	&	"1000"	&	"1110", -- Average = -2
	"0000"	&	"0000"	&	"0000"	&	"1001"	&	"1110", -- Average = -2
	"0000"	&	"0000"	&	"0000"	&	"0000"	&	"0000", -- Average = 0
	"0000"	&	"0000"	&	"0000"	&	"0001"	&	"0000", -- Average = 0
	"0000"	&	"0000"	&	"0000"	&	"0111"	&	"0010", -- Average = 2
	"0000"	&	"0000"	&	"0001"	&	"1000"	&	"1110", -- Average = -2
	"0000"	&	"0000"	&	"0001"	&	"1001"	&	"1110", -- Average = -2
	"0000"	&	"0000"	&	"0001"	&	"0000"	&	"0000", -- Average = 0
	"0000"	&	"0000"	&	"0001"	&	"0001"	&	"0001", -- Average = 1
	"0000"	&	"0000"	&	"0001"	&	"0111"	&	"0010", -- Average = 2
	"0000"	&	"0000"	&	"0111"	&	"1000"	&	"0000", -- Average = 0
	"0000"	&	"0000"	&	"0111"	&	"1001"	&	"0000", -- Average = 0
	"0000"	&	"0000"	&	"0111"	&	"0000"	&	"0010", -- Average = 2
	"0000"	&	"0000"	&	"0111"	&	"0001"	&	"0010", -- Average = 2
	"0000"	&	"0000"	&	"0111"	&	"0111"	&	"0100", -- Average = 4
	"0000"	&	"0001"	&	"1000"	&	"1000"	&	"1100", -- Average = -4
	"0000"	&	"0001"	&	"1000"	&	"1001"	&	"1100", -- Average = -4
	"0000"	&	"0001"	&	"1000"	&	"0000"	&	"1110", -- Average = -2
	"0000"	&	"0001"	&	"1000"	&	"0001"	&	"1110", -- Average = -2
	"0000"	&	"0001"	&	"1000"	&	"0111"	&	"0000", -- Average = 0
	"0000"	&	"0001"	&	"1001"	&	"1000"	&	"1100", -- Average = -4
	"0000"	&	"0001"	&	"1001"	&	"1001"	&	"1101", -- Average = -3
	"0000"	&	"0001"	&	"1001"	&	"0000"	&	"1110", -- Average = -2
	"0000"	&	"0001"	&	"1001"	&	"0001"	&	"1111", -- Average = -1
	"0000"	&	"0001"	&	"1001"	&	"0111"	&	"0000", -- Average = 0
	"0000"	&	"0001"	&	"0000"	&	"1000"	&	"1110", -- Average = -2
	"0000"	&	"0001"	&	"0000"	&	"1001"	&	"1110", -- Average = -2
	"0000"	&	"0001"	&	"0000"	&	"0000"	&	"0000", -- Average = 0
	"0000"	&	"0001"	&	"0000"	&	"0001"	&	"0001", -- Average = 1
	"0000"	&	"0001"	&	"0000"	&	"0111"	&	"0010", -- Average = 2
	"0000"	&	"0001"	&	"0001"	&	"1000"	&	"1110", -- Average = -2
	"0000"	&	"0001"	&	"0001"	&	"1001"	&	"1111", -- Average = -1
	"0000"	&	"0001"	&	"0001"	&	"0000"	&	"0001", -- Average = 1
	"0000"	&	"0001"	&	"0001"	&	"0001"	&	"0001", -- Average = 1
	"0000"	&	"0001"	&	"0001"	&	"0111"	&	"0010", -- Average = 2
	"0000"	&	"0001"	&	"0111"	&	"1000"	&	"0000", -- Average = 0
	"0000"	&	"0001"	&	"0111"	&	"1001"	&	"0000", -- Average = 0
	"0000"	&	"0001"	&	"0111"	&	"0000"	&	"0010", -- Average = 2
	"0000"	&	"0001"	&	"0111"	&	"0001"	&	"0010", -- Average = 2
	"0000"	&	"0001"	&	"0111"	&	"0111"	&	"0100", -- Average = 4
	"0000"	&	"0111"	&	"1000"	&	"1000"	&	"1110", -- Average = -2
	"0000"	&	"0111"	&	"1000"	&	"1001"	&	"1110", -- Average = -2
	"0000"	&	"0111"	&	"1000"	&	"0000"	&	"0000", -- Average = 0
	"0000"	&	"0111"	&	"1000"	&	"0001"	&	"0000", -- Average = 0
	"0000"	&	"0111"	&	"1000"	&	"0111"	&	"0010", -- Average = 2
	"0000"	&	"0111"	&	"1001"	&	"1000"	&	"1110", -- Average = -2
	"0000"	&	"0111"	&	"1001"	&	"1001"	&	"1110", -- Average = -2
	"0000"	&	"0111"	&	"1001"	&	"0000"	&	"0000", -- Average = 0
	"0000"	&	"0111"	&	"1001"	&	"0001"	&	"0000", -- Average = 0
	"0000"	&	"0111"	&	"1001"	&	"0111"	&	"0010", -- Average = 2
	"0000"	&	"0111"	&	"0000"	&	"1000"	&	"0000", -- Average = 0
	"0000"	&	"0111"	&	"0000"	&	"1001"	&	"0000", -- Average = 0
	"0000"	&	"0111"	&	"0000"	&	"0000"	&	"0010", -- Average = 2
	"0000"	&	"0111"	&	"0000"	&	"0001"	&	"0010", -- Average = 2
	"0000"	&	"0111"	&	"0000"	&	"0111"	&	"0100", -- Average = 4
	"0000"	&	"0111"	&	"0001"	&	"1000"	&	"0000", -- Average = 0
	"0000"	&	"0111"	&	"0001"	&	"1001"	&	"0000", -- Average = 0
	"0000"	&	"0111"	&	"0001"	&	"0000"	&	"0010", -- Average = 2
	"0000"	&	"0111"	&	"0001"	&	"0001"	&	"0010", -- Average = 2
	"0000"	&	"0111"	&	"0001"	&	"0111"	&	"0100", -- Average = 4
	"0000"	&	"0111"	&	"0111"	&	"1000"	&	"0010", -- Average = 2
	"0000"	&	"0111"	&	"0111"	&	"1001"	&	"0010", -- Average = 2
	"0000"	&	"0111"	&	"0111"	&	"0000"	&	"0100", -- Average = 4
	"0000"	&	"0111"	&	"0111"	&	"0001"	&	"0100", -- Average = 4
	"0000"	&	"0111"	&	"0111"	&	"0111"	&	"0101", -- Average = 5
	"0001"	&	"1000"	&	"1000"	&	"1000"	&	"1010", -- Average = -6
	"0001"	&	"1000"	&	"1000"	&	"1001"	&	"1010", -- Average = -6
	"0001"	&	"1000"	&	"1000"	&	"0000"	&	"1100", -- Average = -4
	"0001"	&	"1000"	&	"1000"	&	"0001"	&	"1100", -- Average = -4
	"0001"	&	"1000"	&	"1000"	&	"0111"	&	"1110", -- Average = -2
	"0001"	&	"1000"	&	"1001"	&	"1000"	&	"1010", -- Average = -6
	"0001"	&	"1000"	&	"1001"	&	"1001"	&	"1011", -- Average = -5
	"0001"	&	"1000"	&	"1001"	&	"0000"	&	"1100", -- Average = -4
	"0001"	&	"1000"	&	"1001"	&	"0001"	&	"1101", -- Average = -3
	"0001"	&	"1000"	&	"1001"	&	"0111"	&	"1110", -- Average = -2
	"0001"	&	"1000"	&	"0000"	&	"1000"	&	"1100", -- Average = -4
	"0001"	&	"1000"	&	"0000"	&	"1001"	&	"1100", -- Average = -4
	"0001"	&	"1000"	&	"0000"	&	"0000"	&	"1110", -- Average = -2
	"0001"	&	"1000"	&	"0000"	&	"0001"	&	"1110", -- Average = -2
	"0001"	&	"1000"	&	"0000"	&	"0111"	&	"0000", -- Average = 0
	"0001"	&	"1000"	&	"0001"	&	"1000"	&	"1100", -- Average = -4
	"0001"	&	"1000"	&	"0001"	&	"1001"	&	"1101", -- Average = -3
	"0001"	&	"1000"	&	"0001"	&	"0000"	&	"1110", -- Average = -2
	"0001"	&	"1000"	&	"0001"	&	"0001"	&	"1111", -- Average = -1
	"0001"	&	"1000"	&	"0001"	&	"0111"	&	"0000", -- Average = 0
	"0001"	&	"1000"	&	"0111"	&	"1000"	&	"1110", -- Average = -2
	"0001"	&	"1000"	&	"0111"	&	"1001"	&	"1110", -- Average = -2
	"0001"	&	"1000"	&	"0111"	&	"0000"	&	"0000", -- Average = 0
	"0001"	&	"1000"	&	"0111"	&	"0001"	&	"0000", -- Average = 0
	"0001"	&	"1000"	&	"0111"	&	"0111"	&	"0010", -- Average = 2
	"0001"	&	"1001"	&	"1000"	&	"1000"	&	"1010", -- Average = -6
	"0001"	&	"1001"	&	"1000"	&	"1001"	&	"1011", -- Average = -5
	"0001"	&	"1001"	&	"1000"	&	"0000"	&	"1100", -- Average = -4
	"0001"	&	"1001"	&	"1000"	&	"0001"	&	"1101", -- Average = -3
	"0001"	&	"1001"	&	"1000"	&	"0111"	&	"1110", -- Average = -2
	"0001"	&	"1001"	&	"1001"	&	"1000"	&	"1011", -- Average = -5
	"0001"	&	"1001"	&	"1001"	&	"1001"	&	"1011", -- Average = -5
	"0001"	&	"1001"	&	"1001"	&	"0000"	&	"1101", -- Average = -3
	"0001"	&	"1001"	&	"1001"	&	"0001"	&	"1101", -- Average = -3
	"0001"	&	"1001"	&	"1001"	&	"0111"	&	"1110", -- Average = -2
	"0001"	&	"1001"	&	"0000"	&	"1000"	&	"1100", -- Average = -4
	"0001"	&	"1001"	&	"0000"	&	"1001"	&	"1101", -- Average = -3
	"0001"	&	"1001"	&	"0000"	&	"0000"	&	"1110", -- Average = -2
	"0001"	&	"1001"	&	"0000"	&	"0001"	&	"1111", -- Average = -1
	"0001"	&	"1001"	&	"0000"	&	"0111"	&	"0000", -- Average = 0
	"0001"	&	"1001"	&	"0001"	&	"1000"	&	"1101", -- Average = -3
	"0001"	&	"1001"	&	"0001"	&	"1001"	&	"1101", -- Average = -3
	"0001"	&	"1001"	&	"0001"	&	"0000"	&	"1111", -- Average = -1
	"0001"	&	"1001"	&	"0001"	&	"0001"	&	"1111", -- Average = -1
	"0001"	&	"1001"	&	"0001"	&	"0111"	&	"0001", -- Average = 1
	"0001"	&	"1001"	&	"0111"	&	"1000"	&	"1110", -- Average = -2
	"0001"	&	"1001"	&	"0111"	&	"1001"	&	"1110", -- Average = -2
	"0001"	&	"1001"	&	"0111"	&	"0000"	&	"0000", -- Average = 0
	"0001"	&	"1001"	&	"0111"	&	"0001"	&	"0001", -- Average = 1
	"0001"	&	"1001"	&	"0111"	&	"0111"	&	"0010", -- Average = 2
	"0001"	&	"0000"	&	"1000"	&	"1000"	&	"1100", -- Average = -4
	"0001"	&	"0000"	&	"1000"	&	"1001"	&	"1100", -- Average = -4
	"0001"	&	"0000"	&	"1000"	&	"0000"	&	"1110", -- Average = -2
	"0001"	&	"0000"	&	"1000"	&	"0001"	&	"1110", -- Average = -2
	"0001"	&	"0000"	&	"1000"	&	"0111"	&	"0000", -- Average = 0
	"0001"	&	"0000"	&	"1001"	&	"1000"	&	"1100", -- Average = -4
	"0001"	&	"0000"	&	"1001"	&	"1001"	&	"1101", -- Average = -3
	"0001"	&	"0000"	&	"1001"	&	"0000"	&	"1110", -- Average = -2
	"0001"	&	"0000"	&	"1001"	&	"0001"	&	"1111", -- Average = -1
	"0001"	&	"0000"	&	"1001"	&	"0111"	&	"0000", -- Average = 0
	"0001"	&	"0000"	&	"0000"	&	"1000"	&	"1110", -- Average = -2
	"0001"	&	"0000"	&	"0000"	&	"1001"	&	"1110", -- Average = -2
	"0001"	&	"0000"	&	"0000"	&	"0000"	&	"0000", -- Average = 0
	"0001"	&	"0000"	&	"0000"	&	"0001"	&	"0001", -- Average = 1
	"0001"	&	"0000"	&	"0000"	&	"0111"	&	"0010", -- Average = 2
	"0001"	&	"0000"	&	"0001"	&	"1000"	&	"1110", -- Average = -2
	"0001"	&	"0000"	&	"0001"	&	"1001"	&	"1111", -- Average = -1
	"0001"	&	"0000"	&	"0001"	&	"0000"	&	"0001", -- Average = 1
	"0001"	&	"0000"	&	"0001"	&	"0001"	&	"0001", -- Average = 1
	"0001"	&	"0000"	&	"0001"	&	"0111"	&	"0010", -- Average = 2
	"0001"	&	"0000"	&	"0111"	&	"1000"	&	"0000", -- Average = 0
	"0001"	&	"0000"	&	"0111"	&	"1001"	&	"0000", -- Average = 0
	"0001"	&	"0000"	&	"0111"	&	"0000"	&	"0010", -- Average = 2
	"0001"	&	"0000"	&	"0111"	&	"0001"	&	"0010", -- Average = 2
	"0001"	&	"0000"	&	"0111"	&	"0111"	&	"0100", -- Average = 4
	"0001"	&	"0001"	&	"1000"	&	"1000"	&	"1100", -- Average = -4
	"0001"	&	"0001"	&	"1000"	&	"1001"	&	"1101", -- Average = -3
	"0001"	&	"0001"	&	"1000"	&	"0000"	&	"1110", -- Average = -2
	"0001"	&	"0001"	&	"1000"	&	"0001"	&	"1111", -- Average = -1
	"0001"	&	"0001"	&	"1000"	&	"0111"	&	"0000", -- Average = 0
	"0001"	&	"0001"	&	"1001"	&	"1000"	&	"1101", -- Average = -3
	"0001"	&	"0001"	&	"1001"	&	"1001"	&	"1101", -- Average = -3
	"0001"	&	"0001"	&	"1001"	&	"0000"	&	"1111", -- Average = -1
	"0001"	&	"0001"	&	"1001"	&	"0001"	&	"1111", -- Average = -1
	"0001"	&	"0001"	&	"1001"	&	"0111"	&	"0001", -- Average = 1
	"0001"	&	"0001"	&	"0000"	&	"1000"	&	"1110", -- Average = -2
	"0001"	&	"0001"	&	"0000"	&	"1001"	&	"1111", -- Average = -1
	"0001"	&	"0001"	&	"0000"	&	"0000"	&	"0001", -- Average = 1
	"0001"	&	"0001"	&	"0000"	&	"0001"	&	"0001", -- Average = 1
	"0001"	&	"0001"	&	"0000"	&	"0111"	&	"0010", -- Average = 2
	"0001"	&	"0001"	&	"0001"	&	"1000"	&	"1111", -- Average = -1
	"0001"	&	"0001"	&	"0001"	&	"1001"	&	"1111", -- Average = -1
	"0001"	&	"0001"	&	"0001"	&	"0000"	&	"0001", -- Average = 1
	"0001"	&	"0001"	&	"0001"	&	"0001"	&	"0001", -- Average = 1
	"0001"	&	"0001"	&	"0001"	&	"0111"	&	"0011", -- Average = 3
	"0001"	&	"0001"	&	"0111"	&	"1000"	&	"0000", -- Average = 0
	"0001"	&	"0001"	&	"0111"	&	"1001"	&	"0001", -- Average = 1
	"0001"	&	"0001"	&	"0111"	&	"0000"	&	"0010", -- Average = 2
	"0001"	&	"0001"	&	"0111"	&	"0001"	&	"0011", -- Average = 3
	"0001"	&	"0001"	&	"0111"	&	"0111"	&	"0100", -- Average = 4
	"0001"	&	"0111"	&	"1000"	&	"1000"	&	"1110", -- Average = -2
	"0001"	&	"0111"	&	"1000"	&	"1001"	&	"1110", -- Average = -2
	"0001"	&	"0111"	&	"1000"	&	"0000"	&	"0000", -- Average = 0
	"0001"	&	"0111"	&	"1000"	&	"0001"	&	"0000", -- Average = 0
	"0001"	&	"0111"	&	"1000"	&	"0111"	&	"0010", -- Average = 2
	"0001"	&	"0111"	&	"1001"	&	"1000"	&	"1110", -- Average = -2
	"0001"	&	"0111"	&	"1001"	&	"1001"	&	"1110", -- Average = -2
	"0001"	&	"0111"	&	"1001"	&	"0000"	&	"0000", -- Average = 0
	"0001"	&	"0111"	&	"1001"	&	"0001"	&	"0001", -- Average = 1
	"0001"	&	"0111"	&	"1001"	&	"0111"	&	"0010", -- Average = 2
	"0001"	&	"0111"	&	"0000"	&	"1000"	&	"0000", -- Average = 0
	"0001"	&	"0111"	&	"0000"	&	"1001"	&	"0000", -- Average = 0
	"0001"	&	"0111"	&	"0000"	&	"0000"	&	"0010", -- Average = 2
	"0001"	&	"0111"	&	"0000"	&	"0001"	&	"0010", -- Average = 2
	"0001"	&	"0111"	&	"0000"	&	"0111"	&	"0100", -- Average = 4
	"0001"	&	"0111"	&	"0001"	&	"1000"	&	"0000", -- Average = 0
	"0001"	&	"0111"	&	"0001"	&	"1001"	&	"0001", -- Average = 1
	"0001"	&	"0111"	&	"0001"	&	"0000"	&	"0010", -- Average = 2
	"0001"	&	"0111"	&	"0001"	&	"0001"	&	"0011", -- Average = 3
	"0001"	&	"0111"	&	"0001"	&	"0111"	&	"0100", -- Average = 4
	"0001"	&	"0111"	&	"0111"	&	"1000"	&	"0010", -- Average = 2
	"0001"	&	"0111"	&	"0111"	&	"1001"	&	"0010", -- Average = 2
	"0001"	&	"0111"	&	"0111"	&	"0000"	&	"0100", -- Average = 4
	"0001"	&	"0111"	&	"0111"	&	"0001"	&	"0100", -- Average = 4
	"0001"	&	"0111"	&	"0111"	&	"0111"	&	"0110", -- Average = 6
	"0111"	&	"1000"	&	"1000"	&	"1000"	&	"1100", -- Average = -4
	"0111"	&	"1000"	&	"1000"	&	"1001"	&	"1100", -- Average = -4
	"0111"	&	"1000"	&	"1000"	&	"0000"	&	"1110", -- Average = -2
	"0111"	&	"1000"	&	"1000"	&	"0001"	&	"1110", -- Average = -2
	"0111"	&	"1000"	&	"1000"	&	"0111"	&	"1111", -- Average = -1
	"0111"	&	"1000"	&	"1001"	&	"1000"	&	"1100", -- Average = -4
	"0111"	&	"1000"	&	"1001"	&	"1001"	&	"1100", -- Average = -4
	"0111"	&	"1000"	&	"1001"	&	"0000"	&	"1110", -- Average = -2
	"0111"	&	"1000"	&	"1001"	&	"0001"	&	"1110", -- Average = -2
	"0111"	&	"1000"	&	"1001"	&	"0111"	&	"0000", -- Average = 0
	"0111"	&	"1000"	&	"0000"	&	"1000"	&	"1110", -- Average = -2
	"0111"	&	"1000"	&	"0000"	&	"1001"	&	"1110", -- Average = -2
	"0111"	&	"1000"	&	"0000"	&	"0000"	&	"0000", -- Average = 0
	"0111"	&	"1000"	&	"0000"	&	"0001"	&	"0000", -- Average = 0
	"0111"	&	"1000"	&	"0000"	&	"0111"	&	"0010", -- Average = 2
	"0111"	&	"1000"	&	"0001"	&	"1000"	&	"1110", -- Average = -2
	"0111"	&	"1000"	&	"0001"	&	"1001"	&	"1110", -- Average = -2
	"0111"	&	"1000"	&	"0001"	&	"0000"	&	"0000", -- Average = 0
	"0111"	&	"1000"	&	"0001"	&	"0001"	&	"0000", -- Average = 0
	"0111"	&	"1000"	&	"0001"	&	"0111"	&	"0010", -- Average = 2
	"0111"	&	"1000"	&	"0111"	&	"1000"	&	"1111", -- Average = -1
	"0111"	&	"1000"	&	"0111"	&	"1001"	&	"0000", -- Average = 0
	"0111"	&	"1000"	&	"0111"	&	"0000"	&	"0010", -- Average = 2
	"0111"	&	"1000"	&	"0111"	&	"0001"	&	"0010", -- Average = 2
	"0111"	&	"1000"	&	"0111"	&	"0111"	&	"0011", -- Average = 3
	"0111"	&	"1001"	&	"1000"	&	"1000"	&	"1100", -- Average = -4
	"0111"	&	"1001"	&	"1000"	&	"1001"	&	"1100", -- Average = -4
	"0111"	&	"1001"	&	"1000"	&	"0000"	&	"1110", -- Average = -2
	"0111"	&	"1001"	&	"1000"	&	"0001"	&	"1110", -- Average = -2
	"0111"	&	"1001"	&	"1000"	&	"0111"	&	"0000", -- Average = 0
	"0111"	&	"1001"	&	"1001"	&	"1000"	&	"1100", -- Average = -4
	"0111"	&	"1001"	&	"1001"	&	"1001"	&	"1100", -- Average = -4
	"0111"	&	"1001"	&	"1001"	&	"0000"	&	"1110", -- Average = -2
	"0111"	&	"1001"	&	"1001"	&	"0001"	&	"1110", -- Average = -2
	"0111"	&	"1001"	&	"1001"	&	"0111"	&	"0000", -- Average = 0
	"0111"	&	"1001"	&	"0000"	&	"1000"	&	"1110", -- Average = -2
	"0111"	&	"1001"	&	"0000"	&	"1001"	&	"1110", -- Average = -2
	"0111"	&	"1001"	&	"0000"	&	"0000"	&	"0000", -- Average = 0
	"0111"	&	"1001"	&	"0000"	&	"0001"	&	"0000", -- Average = 0
	"0111"	&	"1001"	&	"0000"	&	"0111"	&	"0010", -- Average = 2
	"0111"	&	"1001"	&	"0001"	&	"1000"	&	"1110", -- Average = -2
	"0111"	&	"1001"	&	"0001"	&	"1001"	&	"1110", -- Average = -2
	"0111"	&	"1001"	&	"0001"	&	"0000"	&	"0000", -- Average = 0
	"0111"	&	"1001"	&	"0001"	&	"0001"	&	"0001", -- Average = 1
	"0111"	&	"1001"	&	"0001"	&	"0111"	&	"0010", -- Average = 2
	"0111"	&	"1001"	&	"0111"	&	"1000"	&	"0000", -- Average = 0
	"0111"	&	"1001"	&	"0111"	&	"1001"	&	"0000", -- Average = 0
	"0111"	&	"1001"	&	"0111"	&	"0000"	&	"0010", -- Average = 2
	"0111"	&	"1001"	&	"0111"	&	"0001"	&	"0010", -- Average = 2
	"0111"	&	"1001"	&	"0111"	&	"0111"	&	"0100", -- Average = 4
	"0111"	&	"0000"	&	"1000"	&	"1000"	&	"1110", -- Average = -2
	"0111"	&	"0000"	&	"1000"	&	"1001"	&	"1110", -- Average = -2
	"0111"	&	"0000"	&	"1000"	&	"0000"	&	"0000", -- Average = 0
	"0111"	&	"0000"	&	"1000"	&	"0001"	&	"0000", -- Average = 0
	"0111"	&	"0000"	&	"1000"	&	"0111"	&	"0010", -- Average = 2
	"0111"	&	"0000"	&	"1001"	&	"1000"	&	"1110", -- Average = -2
	"0111"	&	"0000"	&	"1001"	&	"1001"	&	"1110", -- Average = -2
	"0111"	&	"0000"	&	"1001"	&	"0000"	&	"0000", -- Average = 0
	"0111"	&	"0000"	&	"1001"	&	"0001"	&	"0000", -- Average = 0
	"0111"	&	"0000"	&	"1001"	&	"0111"	&	"0010", -- Average = 2
	"0111"	&	"0000"	&	"0000"	&	"1000"	&	"0000", -- Average = 0
	"0111"	&	"0000"	&	"0000"	&	"1001"	&	"0000", -- Average = 0
	"0111"	&	"0000"	&	"0000"	&	"0000"	&	"0010", -- Average = 2
	"0111"	&	"0000"	&	"0000"	&	"0001"	&	"0010", -- Average = 2
	"0111"	&	"0000"	&	"0000"	&	"0111"	&	"0100", -- Average = 4
	"0111"	&	"0000"	&	"0001"	&	"1000"	&	"0000", -- Average = 0
	"0111"	&	"0000"	&	"0001"	&	"1001"	&	"0000", -- Average = 0
	"0111"	&	"0000"	&	"0001"	&	"0000"	&	"0010", -- Average = 2
	"0111"	&	"0000"	&	"0001"	&	"0001"	&	"0010", -- Average = 2
	"0111"	&	"0000"	&	"0001"	&	"0111"	&	"0100", -- Average = 4
	"0111"	&	"0000"	&	"0111"	&	"1000"	&	"0010", -- Average = 2
	"0111"	&	"0000"	&	"0111"	&	"1001"	&	"0010", -- Average = 2
	"0111"	&	"0000"	&	"0111"	&	"0000"	&	"0100", -- Average = 4
	"0111"	&	"0000"	&	"0111"	&	"0001"	&	"0100", -- Average = 4
	"0111"	&	"0000"	&	"0111"	&	"0111"	&	"0101", -- Average = 5
	"0111"	&	"0001"	&	"1000"	&	"1000"	&	"1110", -- Average = -2
	"0111"	&	"0001"	&	"1000"	&	"1001"	&	"1110", -- Average = -2
	"0111"	&	"0001"	&	"1000"	&	"0000"	&	"0000", -- Average = 0
	"0111"	&	"0001"	&	"1000"	&	"0001"	&	"0000", -- Average = 0
	"0111"	&	"0001"	&	"1000"	&	"0111"	&	"0010", -- Average = 2
	"0111"	&	"0001"	&	"1001"	&	"1000"	&	"1110", -- Average = -2
	"0111"	&	"0001"	&	"1001"	&	"1001"	&	"1110", -- Average = -2
	"0111"	&	"0001"	&	"1001"	&	"0000"	&	"0000", -- Average = 0
	"0111"	&	"0001"	&	"1001"	&	"0001"	&	"0001", -- Average = 1
	"0111"	&	"0001"	&	"1001"	&	"0111"	&	"0010", -- Average = 2
	"0111"	&	"0001"	&	"0000"	&	"1000"	&	"0000", -- Average = 0
	"0111"	&	"0001"	&	"0000"	&	"1001"	&	"0000", -- Average = 0
	"0111"	&	"0001"	&	"0000"	&	"0000"	&	"0010", -- Average = 2
	"0111"	&	"0001"	&	"0000"	&	"0001"	&	"0010", -- Average = 2
	"0111"	&	"0001"	&	"0000"	&	"0111"	&	"0100", -- Average = 4
	"0111"	&	"0001"	&	"0001"	&	"1000"	&	"0000", -- Average = 0
	"0111"	&	"0001"	&	"0001"	&	"1001"	&	"0001", -- Average = 1
	"0111"	&	"0001"	&	"0001"	&	"0000"	&	"0010", -- Average = 2
	"0111"	&	"0001"	&	"0001"	&	"0001"	&	"0011", -- Average = 3
	"0111"	&	"0001"	&	"0001"	&	"0111"	&	"0100", -- Average = 4
	"0111"	&	"0001"	&	"0111"	&	"1000"	&	"0010", -- Average = 2
	"0111"	&	"0001"	&	"0111"	&	"1001"	&	"0010", -- Average = 2
	"0111"	&	"0001"	&	"0111"	&	"0000"	&	"0100", -- Average = 4
	"0111"	&	"0001"	&	"0111"	&	"0001"	&	"0100", -- Average = 4
	"0111"	&	"0001"	&	"0111"	&	"0111"	&	"0110", -- Average = 6
	"0111"	&	"0111"	&	"1000"	&	"1000"	&	"1111", -- Average = -1
	"0111"	&	"0111"	&	"1000"	&	"1001"	&	"0000", -- Average = 0
	"0111"	&	"0111"	&	"1000"	&	"0000"	&	"0010", -- Average = 2
	"0111"	&	"0111"	&	"1000"	&	"0001"	&	"0010", -- Average = 2
	"0111"	&	"0111"	&	"1000"	&	"0111"	&	"0011", -- Average = 3
	"0111"	&	"0111"	&	"1001"	&	"1000"	&	"0000", -- Average = 0
	"0111"	&	"0111"	&	"1001"	&	"1001"	&	"0000", -- Average = 0
	"0111"	&	"0111"	&	"1001"	&	"0000"	&	"0010", -- Average = 2
	"0111"	&	"0111"	&	"1001"	&	"0001"	&	"0010", -- Average = 2
	"0111"	&	"0111"	&	"1001"	&	"0111"	&	"0100", -- Average = 4
	"0111"	&	"0111"	&	"0000"	&	"1000"	&	"0010", -- Average = 2
	"0111"	&	"0111"	&	"0000"	&	"1001"	&	"0010", -- Average = 2
	"0111"	&	"0111"	&	"0000"	&	"0000"	&	"0100", -- Average = 4
	"0111"	&	"0111"	&	"0000"	&	"0001"	&	"0100", -- Average = 4
	"0111"	&	"0111"	&	"0000"	&	"0111"	&	"0101", -- Average = 5
	"0111"	&	"0111"	&	"0001"	&	"1000"	&	"0010", -- Average = 2
	"0111"	&	"0111"	&	"0001"	&	"1001"	&	"0010", -- Average = 2
	"0111"	&	"0111"	&	"0001"	&	"0000"	&	"0100", -- Average = 4
	"0111"	&	"0111"	&	"0001"	&	"0001"	&	"0100", -- Average = 4
	"0111"	&	"0111"	&	"0001"	&	"0111"	&	"0110", -- Average = 6
	"0111"	&	"0111"	&	"0111"	&	"1000"	&	"0011", -- Average = 3
	"0111"	&	"0111"	&	"0111"	&	"1001"	&	"0100", -- Average = 4
	"0111"	&	"0111"	&	"0111"	&	"0000"	&	"0101", -- Average = 5
	"0111"	&	"0111"	&	"0111"	&	"0001"	&	"0110", -- Average = 6
	"0111"	&	"0111"	&	"0111"	&	"0111"	&	"0111" -- Average = 7
	);
 
BEGIN
 
 
	-- Instantiate the Unit Under Test (UUT)
   uut: FindAverage_4bit PORT MAP (
          A => A,
          B => B,
          C => C,
          D => D,
          AVERAGE => AVERAGE
        );

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      for i in test_vector'Range loop
			
			A <= test_vector(i)(19 downto 16);
			B <= test_vector(i)(15 downto 12);
			C <= test_vector(i)(11 downto 8);
			D <= test_vector(i)(7 downto 4);
			
			wait for 20 ns;
			
			assert ( AVERAGE = test_vector(i)(3 downto 0))
			report "***** Test failed. *****"
         severity Failure;
			
		end loop;
      
		
		      -- All tests are successful if we get this far
      report "***** All tests completed successfully. *****";
      wait;
   end process;

END;
