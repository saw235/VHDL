----------------------------------------------------------------------------
-- Entity:        CompareEQU_4bit_tb
-- Written By:    Saw Xue Zheng
-- Date Created:  9/11/2016
-- Description:   Testbench for CompareEQU_4bit
--
-- Revision History (date, initials, description):
-- 	11 Sept 16, xps5001, file created.

-- Dependencies:
--		CompareEQU_4bit
----------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
 
ENTITY CompareEQU_4bit_tb IS
END CompareEQU_4bit_tb;
 
ARCHITECTURE behavior OF CompareEQU_4bit_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT CompareEQU_4bit
    PORT(
         A   : IN  std_logic_vector(3 downto 0);
         B   : IN  std_logic_vector(3 downto 0);
         EQU : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic_vector(3 downto 0) := (others => '0');
   signal B : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal EQU : std_logic;

   type test_vector_type is array (0 to 255) of STD_LOGIC_VECTOR (8 downto 0);
	constant test_vector : test_vector_type := (
	 --A          B          EQU
	"0000"	&	"0000"	&	"1",
	"0000"	&	"0001"	&	"0",
	"0000"	&	"0010"	&	"0",
	"0000"	&	"0011"	&	"0",
	"0000"	&	"0100"	&	"0",
	"0000"	&	"0101"	&	"0",
	"0000"	&	"0110"	&	"0",
	"0000"	&	"0111"	&	"0",
	"0000"	&	"1000"	&	"0",
	"0000"	&	"1001"	&	"0",
	"0000"	&	"1010"	&	"0",
	"0000"	&	"1011"	&	"0",
	"0000"	&	"1100"	&	"0",
	"0000"	&	"1101"	&	"0",
	"0000"	&	"1110"	&	"0",
	"0000"	&	"1111"	&	"0",
	"0001"	&	"0000"	&	"0",
	"0001"	&	"0001"	&	"1",
	"0001"	&	"0010"	&	"0",
	"0001"	&	"0011"	&	"0",
	"0001"	&	"0100"	&	"0",
	"0001"	&	"0101"	&	"0",
	"0001"	&	"0110"	&	"0",
	"0001"	&	"0111"	&	"0",
	"0001"	&	"1000"	&	"0",
	"0001"	&	"1001"	&	"0",
	"0001"	&	"1010"	&	"0",
	"0001"	&	"1011"	&	"0",
	"0001"	&	"1100"	&	"0",
	"0001"	&	"1101"	&	"0",
	"0001"	&	"1110"	&	"0",
	"0001"	&	"1111"	&	"0",
	"0010"	&	"0000"	&	"0",
	"0010"	&	"0001"	&	"0",
	"0010"	&	"0010"	&	"1",
	"0010"	&	"0011"	&	"0",
	"0010"	&	"0100"	&	"0",
	"0010"	&	"0101"	&	"0",
	"0010"	&	"0110"	&	"0",
	"0010"	&	"0111"	&	"0",
	"0010"	&	"1000"	&	"0",
	"0010"	&	"1001"	&	"0",
	"0010"	&	"1010"	&	"0",
	"0010"	&	"1011"	&	"0",
	"0010"	&	"1100"	&	"0",
	"0010"	&	"1101"	&	"0",
	"0010"	&	"1110"	&	"0",
	"0010"	&	"1111"	&	"0",
	"0011"	&	"0000"	&	"0",
	"0011"	&	"0001"	&	"0",
	"0011"	&	"0010"	&	"0",
	"0011"	&	"0011"	&	"1",
	"0011"	&	"0100"	&	"0",
	"0011"	&	"0101"	&	"0",
	"0011"	&	"0110"	&	"0",
	"0011"	&	"0111"	&	"0",
	"0011"	&	"1000"	&	"0",
	"0011"	&	"1001"	&	"0",
	"0011"	&	"1010"	&	"0",
	"0011"	&	"1011"	&	"0",
	"0011"	&	"1100"	&	"0",
	"0011"	&	"1101"	&	"0",
	"0011"	&	"1110"	&	"0",
	"0011"	&	"1111"	&	"0",
	"0100"	&	"0000"	&	"0",
	"0100"	&	"0001"	&	"0",
	"0100"	&	"0010"	&	"0",
	"0100"	&	"0011"	&	"0",
	"0100"	&	"0100"	&	"1",
	"0100"	&	"0101"	&	"0",
	"0100"	&	"0110"	&	"0",
	"0100"	&	"0111"	&	"0",
	"0100"	&	"1000"	&	"0",
	"0100"	&	"1001"	&	"0",
	"0100"	&	"1010"	&	"0",
	"0100"	&	"1011"	&	"0",
	"0100"	&	"1100"	&	"0",
	"0100"	&	"1101"	&	"0",
	"0100"	&	"1110"	&	"0",
	"0100"	&	"1111"	&	"0",
	"0101"	&	"0000"	&	"0",
	"0101"	&	"0001"	&	"0",
	"0101"	&	"0010"	&	"0",
	"0101"	&	"0011"	&	"0",
	"0101"	&	"0100"	&	"0",
	"0101"	&	"0101"	&	"1",
	"0101"	&	"0110"	&	"0",
	"0101"	&	"0111"	&	"0",
	"0101"	&	"1000"	&	"0",
	"0101"	&	"1001"	&	"0",
	"0101"	&	"1010"	&	"0",
	"0101"	&	"1011"	&	"0",
	"0101"	&	"1100"	&	"0",
	"0101"	&	"1101"	&	"0",
	"0101"	&	"1110"	&	"0",
	"0101"	&	"1111"	&	"0",
	"0110"	&	"0000"	&	"0",
	"0110"	&	"0001"	&	"0",
	"0110"	&	"0010"	&	"0",
	"0110"	&	"0011"	&	"0",
	"0110"	&	"0100"	&	"0",
	"0110"	&	"0101"	&	"0",
	"0110"	&	"0110"	&	"1",
	"0110"	&	"0111"	&	"0",
	"0110"	&	"1000"	&	"0",
	"0110"	&	"1001"	&	"0",
	"0110"	&	"1010"	&	"0",
	"0110"	&	"1011"	&	"0",
	"0110"	&	"1100"	&	"0",
	"0110"	&	"1101"	&	"0",
	"0110"	&	"1110"	&	"0",
	"0110"	&	"1111"	&	"0",
	"0111"	&	"0000"	&	"0",
	"0111"	&	"0001"	&	"0",
	"0111"	&	"0010"	&	"0",
	"0111"	&	"0011"	&	"0",
	"0111"	&	"0100"	&	"0",
	"0111"	&	"0101"	&	"0",
	"0111"	&	"0110"	&	"0",
	"0111"	&	"0111"	&	"1",
	"0111"	&	"1000"	&	"0",
	"0111"	&	"1001"	&	"0",
	"0111"	&	"1010"	&	"0",
	"0111"	&	"1011"	&	"0",
	"0111"	&	"1100"	&	"0",
	"0111"	&	"1101"	&	"0",
	"0111"	&	"1110"	&	"0",
	"0111"	&	"1111"	&	"0",
	"1000"	&	"0000"	&	"0",
	"1000"	&	"0001"	&	"0",
	"1000"	&	"0010"	&	"0",
	"1000"	&	"0011"	&	"0",
	"1000"	&	"0100"	&	"0",
	"1000"	&	"0101"	&	"0",
	"1000"	&	"0110"	&	"0",
	"1000"	&	"0111"	&	"0",
	"1000"	&	"1000"	&	"1",
	"1000"	&	"1001"	&	"0",
	"1000"	&	"1010"	&	"0",
	"1000"	&	"1011"	&	"0",
	"1000"	&	"1100"	&	"0",
	"1000"	&	"1101"	&	"0",
	"1000"	&	"1110"	&	"0",
	"1000"	&	"1111"	&	"0",
	"1001"	&	"0000"	&	"0",
	"1001"	&	"0001"	&	"0",
	"1001"	&	"0010"	&	"0",
	"1001"	&	"0011"	&	"0",
	"1001"	&	"0100"	&	"0",
	"1001"	&	"0101"	&	"0",
	"1001"	&	"0110"	&	"0",
	"1001"	&	"0111"	&	"0",
	"1001"	&	"1000"	&	"0",
	"1001"	&	"1001"	&	"1",
	"1001"	&	"1010"	&	"0",
	"1001"	&	"1011"	&	"0",
	"1001"	&	"1100"	&	"0",
	"1001"	&	"1101"	&	"0",
	"1001"	&	"1110"	&	"0",
	"1001"	&	"1111"	&	"0",
	"1010"	&	"0000"	&	"0",
	"1010"	&	"0001"	&	"0",
	"1010"	&	"0010"	&	"0",
	"1010"	&	"0011"	&	"0",
	"1010"	&	"0100"	&	"0",
	"1010"	&	"0101"	&	"0",
	"1010"	&	"0110"	&	"0",
	"1010"	&	"0111"	&	"0",
	"1010"	&	"1000"	&	"0",
	"1010"	&	"1001"	&	"0",
	"1010"	&	"1010"	&	"1",
	"1010"	&	"1011"	&	"0",
	"1010"	&	"1100"	&	"0",
	"1010"	&	"1101"	&	"0",
	"1010"	&	"1110"	&	"0",
	"1010"	&	"1111"	&	"0",
	"1011"	&	"0000"	&	"0",
	"1011"	&	"0001"	&	"0",
	"1011"	&	"0010"	&	"0",
	"1011"	&	"0011"	&	"0",
	"1011"	&	"0100"	&	"0",
	"1011"	&	"0101"	&	"0",
	"1011"	&	"0110"	&	"0",
	"1011"	&	"0111"	&	"0",
	"1011"	&	"1000"	&	"0",
	"1011"	&	"1001"	&	"0",
	"1011"	&	"1010"	&	"0",
	"1011"	&	"1011"	&	"1",
	"1011"	&	"1100"	&	"0",
	"1011"	&	"1101"	&	"0",
	"1011"	&	"1110"	&	"0",
	"1011"	&	"1111"	&	"0",
	"1100"	&	"0000"	&	"0",
	"1100"	&	"0001"	&	"0",
	"1100"	&	"0010"	&	"0",
	"1100"	&	"0011"	&	"0",
	"1100"	&	"0100"	&	"0",
	"1100"	&	"0101"	&	"0",
	"1100"	&	"0110"	&	"0",
	"1100"	&	"0111"	&	"0",
	"1100"	&	"1000"	&	"0",
	"1100"	&	"1001"	&	"0",
	"1100"	&	"1010"	&	"0",
	"1100"	&	"1011"	&	"0",
	"1100"	&	"1100"	&	"1",
	"1100"	&	"1101"	&	"0",
	"1100"	&	"1110"	&	"0",
	"1100"	&	"1111"	&	"0",
	"1101"	&	"0000"	&	"0",
	"1101"	&	"0001"	&	"0",
	"1101"	&	"0010"	&	"0",
	"1101"	&	"0011"	&	"0",
	"1101"	&	"0100"	&	"0",
	"1101"	&	"0101"	&	"0",
	"1101"	&	"0110"	&	"0",
	"1101"	&	"0111"	&	"0",
	"1101"	&	"1000"	&	"0",
	"1101"	&	"1001"	&	"0",
	"1101"	&	"1010"	&	"0",
	"1101"	&	"1011"	&	"0",
	"1101"	&	"1100"	&	"0",
	"1101"	&	"1101"	&	"1",
	"1101"	&	"1110"	&	"0",
	"1101"	&	"1111"	&	"0",
	"1110"	&	"0000"	&	"0",
	"1110"	&	"0001"	&	"0",
	"1110"	&	"0010"	&	"0",
	"1110"	&	"0011"	&	"0",
	"1110"	&	"0100"	&	"0",
	"1110"	&	"0101"	&	"0",
	"1110"	&	"0110"	&	"0",
	"1110"	&	"0111"	&	"0",
	"1110"	&	"1000"	&	"0",
	"1110"	&	"1001"	&	"0",
	"1110"	&	"1010"	&	"0",
	"1110"	&	"1011"	&	"0",
	"1110"	&	"1100"	&	"0",
	"1110"	&	"1101"	&	"0",
	"1110"	&	"1110"	&	"1",
	"1110"	&	"1111"	&	"0",
	"1111"	&	"0000"	&	"0",
	"1111"	&	"0001"	&	"0",
	"1111"	&	"0010"	&	"0",
	"1111"	&	"0011"	&	"0",
	"1111"	&	"0100"	&	"0",
	"1111"	&	"0101"	&	"0",
	"1111"	&	"0110"	&	"0",
	"1111"	&	"0111"	&	"0",
	"1111"	&	"1000"	&	"0",
	"1111"	&	"1001"	&	"0",
	"1111"	&	"1010"	&	"0",
	"1111"	&	"1011"	&	"0",
	"1111"	&	"1100"	&	"0",
	"1111"	&	"1101"	&	"0",
	"1111"	&	"1110"	&	"0",
	"1111"	&	"1111"	&	"1"
	);
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: CompareEQU_4bit PORT MAP (
          A => A,
          B => B,
          EQU => EQU
        );
 

   -- Stimulus process
   stim_proc: process
   begin

      -- hold reset state for 100 ns.
      wait for 100 ns;
		
		-- run through all test vectors
      for i in test_vector'Range loop
      
         -- Assign test inputs
         A <= test_vector(i)(8 downto 5);
         B <= test_vector(i)(4 downto 1);
         -- Compare outputs to expected values
         wait for 2ns;
         assert (EQU = test_vector(i)(0))
            report "***** Test failed. *****"
            severity Failure;
      end loop;
      
      -- All tests are successful if we get this far
      report "***** All tests completed successfully. *****";
      wait;
   end process;

END;
